ENTITY SHIFT_REG IS
	GENERIC(N : INTEGER := 8);
	PORT (
			CLK		: IN BIT;
			DIN		: IN INTEGER;
			DOUT	: OUT INTEGER
	);
END ENTITY SHIFT_REG;

ARCHITECTURE BEHAVIOR OF SHIFT_REG IS
	TYPE INT_ARRAY IS ARRAY (N DOWN TO 0) OF INTEGER;
	SIGNAL	D_REG : INT_ARRAY;
	BEGIN
		PROCESS (CLK) IS
			BEGIN
				IF (CLK'EVENT AND CLK='1') THEN
					D_RED<=DIN & D_REG(N DOWNTO 1);
				END IF;
		END PROCESS;
		DOUT<=D_REG(0);
END ARCHITECTURE BEHAVIOR;

----------------------------------------- TESTBENCH

ENTITY TB IS
GENERIC (N : INTEGER = 4);
END ENTITY TB;

ARCHITECTURE TB OF TB IS
	SIGNAL S_DIN, S_DOUT BIT;
	SIGNAL S_CLK : BIT :='0';
	BEGIN
		DUT:ENTITY SHIFT_REG (BEHAVIOR)
		GENERIC MAP(N)
		PORT MAP(S_CLK,S_DIN,S_DOUT);
		
		S_CLK<=NOT S_CLK AFTER 50 NS;
		
		PROCESS IS
			BEGIN
			S_DIN<=	69,
					90 AFTER 125 NS,
					100 AFTER 225 NS,
					669 AFTER 325 NS,
					789 AFTER 425 NS;
			WAIT FOR 500 NS;
		END PROCESS;
END ARCHITECTURE;