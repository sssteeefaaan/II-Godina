LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;		--TO_INTEGER (UNSIGNED)
--USE IEEE.STD_LOGIC_ARITH.ALL;	--CONV_INTEGER(UNSIGNED)


ENTITY DECODER IS
GENERIC (N: INTEGER:=4);
PORT(
	ENABLE	: IN BIT;
	Xin		: IN STD_LOGIC_VECTOR (N-1 DOWNTO 0);
	Yout	: OUT STD_LOGIC_VECTOR (2**N-1 DOWNTO 0)
);
END ENTITY DECODER;

ARCHITECTURE BEHAVIOR OF DECODER IS
	BEGIN
		PROCESS (ENABLE,Xin)
          VARIABLE ADRESS: INTEGER RANGE 0 TO 2**N-1;
          VARIABLE OUTPUT: STD_LOGIC_VECTOR (2**N-1 DOWNTO 0);
          BEGIN
              OUTPUT:=(OTHERS=>'1');
              IF(ENABLE='1') THEN
                  ADRESS:=TO_INTEGER(UNSIGNED(Xin));
                  OUTPUT(ADRESS):='0';
              END IF;
              Yout<=OUTPUT;
		END PROCESS;
END ARCHITECTURE BEHAVIOR;

----------------------------------------------------  BEZ PROMENLJIVIH

ARCHITECTURE BEHAVIORDIRECT OF DECODER IS
	BEGIN
		PROCESS (ENABLE,Xin)
          BEGIN
              Yout=(OTHERS=>'1');
              IF(ENABLE='1') THEN
                  Yout(TO_INTEGER(UNSIGNED(Xin)))<='0';
              END IF;
		END PROCESS;
END ARCHITECTURE BEHAVIOR;

--------------------------------------------- TESTBENCH

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
--USE IEEE.NUMERIC_STD.ALL; -- NE SMEJU OBA

ENTITY TB IS
GENERIC (N:INTEGER:=4);
END ENTITY TB;

ARCHITECTURE TB OF TB IS
SIGNAL S_ENABLE : BIT;
SIGNAL S_Xin	: STD_LOGIC_VECTOR (N-1 DOWNTO 0);
SIGNAL S_Yout	: STD_LOGIC_VECTOR (2**N-1 DOWNTO 0);

	BEGIN
		DUT: ENTITY DECODER(BEHAVIOR)
		GENERIC MAP(N)
		PORT MAP(S_ENABLE,S_Xin,S_Yout);
		
		TEST: PROCESS IS
			BEGIN
				S_ENABLE<='0', '1' AFTER 10 NS;
				S_Xin<="0000"; -- 0
				WAIT FOR 25 NS;
				S_Xin<="0100"; -- 4
				WAIT FOR 25 NS;
                S_Xin<="1000"; -- 8
				WAIT FOR 25 NS;
				S_Xin<="1100"; -- 12
				WAIT FOR 25 NS;
		END PROCESS TEST;
END ARCHITECTURE TB;